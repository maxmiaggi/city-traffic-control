library verilog;
use verilog.vl_types.all;
entity level1_tb is
end level1_tb;
