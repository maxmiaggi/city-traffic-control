library verilog;
use verilog.vl_types.all;
entity randomtest1_tb is
end randomtest1_tb;
